`timescale 1ns/1ns
module tone_generator (
    input clk,
    input output_enable,
    input [23:0] tone_switch_period,
    input volume,
    output square_wave_out
);
    // TODO(you): Your code here. Remove the following lines once you add your implementation.
    assign square_wave_out = 1'b0;
endmodule
